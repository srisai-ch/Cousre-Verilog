`include "half_adder_gate.v"
`include "full_adder_using_ha.v"
`include "tb_full_adder.v"